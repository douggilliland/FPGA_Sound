-- Middle C sine wave table
-- 50 MHz Clock
-- 8 bit PWM samples
-- Clock prescaler = 4, 12.5 MHz
-- 12.5 MHz / 256 = 48828.125 KHz
-- Middle C is 261.626 Hz

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

ENTITY MiddleCSine8Table IS
	PORT
	(
		address : in std_logic_vector(7 downto 0);
		q : out std_logic_vector(7 downto 0)
	);
END MiddleCSine8Table;

architecture behavior of MiddleCSine8Table is
type romtable is array (0 to 186) of std_logic_vector(7 downto 0);
constant romdata : romtable :=
(
x"7F",
x"83",
x"88",
x"8C",
x"90",
x"94",
x"98",
x"9D",
x"A1",
x"A5",
x"A9",
x"AD",
x"B1",
x"B5",
x"B9",
x"BC",
x"C0",
x"C4",
x"C7",
x"CB",
x"CE",
x"D1",
x"D5",
x"D8",
x"DB",
x"DE",
x"E0",
x"E3",
x"E6",
x"E8",
x"EA",
x"ED",
x"EF",
x"F1",
x"F3",
x"F4",
x"F6",
x"F7",
x"F9",
x"FA",
x"FB",
x"FC",
x"FC",
x"FD",
x"FD",
x"FE",
x"FE",
x"FE",
x"FE",
x"FE",
x"FD",
x"FD",
x"FC",
x"FB",
x"FA",
x"F9",
x"F8",
x"F7",
x"F5",
x"F3",
x"F2",
x"F0",
x"EE",
x"EC",
x"E9",
x"E7",
x"E4",
x"E2",
x"DF",
x"DC",
x"D9",
x"D6",
x"D3",
x"D0",
x"CC",
x"C9",
x"C5",
x"C2",
x"BE",
x"BA",
x"B7",
x"B3",
x"AF",
x"AB",
x"A7",
x"A3",
x"9F",
x"9B",
x"96",
x"92",
x"8E",
x"8A",
x"85",
x"81",
x"7D",
x"79",
x"74",
x"70",
x"6C",
x"68",
x"63",
x"5F",
x"5B",
x"57",
x"53",
x"4F",
x"4B",
x"47",
x"44",
x"40",
x"3C",
x"39",
x"35",
x"32",
x"2E",
x"2B",
x"28",
x"25",
x"22",
x"1F",
x"1C",
x"1A",
x"17",
x"15",
x"12",
x"10",
x"0E",
x"0C",
x"0B",
x"09",
x"07",
x"06",
x"05",
x"04",
x"03",
x"02",
x"01",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"01",
x"02",
x"02",
x"03",
x"04",
x"05",
x"07",
x"08",
x"0A",
x"0B",
x"0D",
x"0F",
x"11",
x"14",
x"16",
x"18",
x"1B",
x"1E",
x"20",
x"23",
x"26",
x"29",
x"2D",
x"30",
x"33",
x"37",
x"3A",
x"3E",
x"42",
x"45",
x"49",
x"4D",
x"51",
x"55",
x"59",
x"5D",
x"61",
x"66",
x"6A",
x"6E",
x"72",
x"76",
x"7B"
);
begin
process (address)
begin
q <= romdata (to_integer(unsigned(address)));
end process;
end behavior;
