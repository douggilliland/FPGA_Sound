-- Middle C sine wave table
-- 50 MHz Clock
-- 8 bit PWM samples
-- 256 samples contain entire sine wave
-- Middle C is 261.626 Hz

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

ENTITY MiddleCSine8Table IS
	PORT
	(
		address : in std_logic_vector(7 downto 0);
		q : out std_logic_vector(7 downto 0)
	);
END MiddleCSine8Table;

architecture behavior of MiddleCSine8Table is
type romtable is array (0 to 255) of std_logic_vector(7 downto 0);
constant romdata : romtable :=
(
x"7F",
x"82",
x"85",
x"88",
x"8B",
x"8F",
x"92",
x"95",
x"98",
x"9B",
x"9E",
x"A1",
x"A4",
x"A7",
x"AA",
x"AD",
x"B0",
x"B2",
x"B5",
x"B8",
x"BB",
x"BE",
x"C0",
x"C3",
x"C6",
x"C8",
x"CB",
x"CD",
x"D0",
x"D2",
x"D4",
x"D7",
x"D9",
x"DB",
x"DD",
x"DF",
x"E1",
x"E3",
x"E5",
x"E7",
x"E9",
x"EA",
x"EC",
x"EE",
x"EF",
x"F0",
x"F2",
x"F3",
x"F4",
x"F5",
x"F7",
x"F8",
x"F9",
x"F9",
x"FA",
x"FB",
x"FC",
x"FC",
x"FD",
x"FD",
x"FD",
x"FE",
x"FE",
x"FE",
x"FE",
x"FE",
x"FE",
x"FE",
x"FD",
x"FD",
x"FD",
x"FC",
x"FC",
x"FB",
x"FA",
x"F9",
x"F9",
x"F8",
x"F7",
x"F5",
x"F4",
x"F3",
x"F2",
x"F0",
x"EF",
x"EE",
x"EC",
x"EA",
x"E9",
x"E7",
x"E5",
x"E3",
x"E1",
x"DF",
x"DD",
x"DB",
x"D9",
x"D7",
x"D4",
x"D2",
x"D0",
x"CD",
x"CB",
x"C8",
x"C6",
x"C3",
x"C0",
x"BE",
x"BB",
x"B8",
x"B5",
x"B2",
x"B0",
x"AD",
x"AA",
x"A7",
x"A4",
x"A1",
x"9E",
x"9B",
x"98",
x"95",
x"92",
x"8F",
x"8B",
x"88",
x"85",
x"82",
x"7F",
x"7C",
x"79",
x"76",
x"73",
x"6F",
x"6C",
x"69",
x"66",
x"63",
x"60",
x"5D",
x"5A",
x"57",
x"54",
x"51",
x"4E",
x"4C",
x"49",
x"46",
x"43",
x"40",
x"3E",
x"3B",
x"38",
x"36",
x"33",
x"31",
x"2E",
x"2C",
x"2A",
x"27",
x"25",
x"23",
x"21",
x"1F",
x"1D",
x"1B",
x"19",
x"17",
x"15",
x"14",
x"12",
x"10",
x"0F",
x"0E",
x"0C",
x"0B",
x"0A",
x"09",
x"07",
x"06",
x"05",
x"05",
x"04",
x"03",
x"02",
x"02",
x"01",
x"01",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"01",
x"01",
x"02",
x"02",
x"03",
x"04",
x"05",
x"05",
x"06",
x"07",
x"09",
x"0A",
x"0B",
x"0C",
x"0E",
x"0F",
x"10",
x"12",
x"14",
x"15",
x"17",
x"19",
x"1B",
x"1D",
x"1F",
x"21",
x"23",
x"25",
x"27",
x"2A",
x"2C",
x"2E",
x"31",
x"33",
x"36",
x"38",
x"3B",
x"3E",
x"40",
x"43",
x"46",
x"49",
x"4C",
x"4E",
x"51",
x"54",
x"57",
x"5A",
x"5D",
x"60",
x"63",
x"66",
x"69",
x"6C",
x"6F",
x"73",
x"76",
x"79",
x"7C"
);
begin
process (address)
begin
q <= romdata (to_integer(unsigned(address)));
end process;
end behavior;
